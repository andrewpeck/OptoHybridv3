----------------------------------------------------------------------------------
-- CMS Muon Endcap
-- GEM Collaboration
-- Optohybrid v3 Firmware -- Clocking
-- A. Peck
----------------------------------------------------------------------------------
-- 2017/07/21 -- Initial port to version 3 electronics
-- 2017/07/22 -- Additional MMCM added to monitor and dejitter the eport clock
-- 2017/08/09 -- 200MHz iodelay refclk added to primary MMCM
-- 2019/05/02 -- Added BUFGCE outputs to disable clocks during MGT init
-- 2019/05/09 -- Cleanup clocking with new gated clocking scheme
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_misc.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.types_pkg.all;
use work.param_pkg.all;
use work.ipbus_pkg.all;
use work.registers.all;

entity clocking is
generic(
    g_ERROR_COUNT_MAX : integer := 5;
    g_DONT_USE_CLOCK_GATING : std_logic := '0'
);
port(

    -- gbt_eclk_p  : in std_logic_vector (1 downto 0);
    -- gbt_eclk_n  : in std_logic_vector (1 downto 0);

    -- programmable frequency/phase deskew clocks
    clock_i_p : in std_logic;
    clock_i_n : in std_logic;

    -- logic clocks
    clk_1x_o: out std_logic;
    clk_2x_o: out std_logic;
    clk_4x_o: out std_logic;
    clk_4x_90_o: out std_logic;
    clk_5x_o: out std_logic;

    clk_1x_gated_o          : out std_logic;
    clk_2x_gated_o          : out std_logic;
    clk_4x_gated_o          : out std_logic;
    clk_4x_90_gated_o       : out std_logic;
    clk_5x_gated_o          : out std_logic;

    -- mmcm locked status monitors
    trigger_mmcm_locked_o   : out std_logic;
    core_mmcm_locked_o   : out std_logic;

    mmcms_locked_o   : out std_logic;

    clock_enable_i  : in std_logic;

    -- ipbus

    ipb_mosi_i : in  ipb_wbus;
    ipb_miso_o : out ipb_rbus;

    ipb_reset_i : in std_logic;

    sump : out std_logic

);
end clocking;


architecture Behavioral of clocking is

    signal mmcm_locked : std_logic_vector(1 downto 0);
    signal mmcm_unlocked : std_logic_vector(1 downto 0);

    signal clock_i : std_logic;
    signal clock   : std_logic;

    ------ Register signals begin (this section is generated by <optohybrid_top>/tools/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_write_arr       : t_std32_array(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_addresses       : t_std32_array(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_defaults        : t_std32_array(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_write_arr_sump  : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0);
    signal regs_read_pulse_arr  : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '0');
    signal regs_write_pulse_arr : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '0');
    signal regs_read_ready_arr  : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '0');
    -- Connect counter signal declarations
    signal cnt_gbt_mmcm_unlocked : std_logic_vector (7 downto 0) := (others => '0');
    signal cnt_logic_mmcm_unlocked : std_logic_vector (7 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------

begin

    clk_1x_o          <= clock;

    mmcm_unlocked <= not mmcm_locked;

    mmcms_locked_o     <= mmcm_locked(0) and mmcm_locked(1);

    trigger_mmcm_locked_o <= mmcm_locked(0);
    core_mmcm_locked_o <= mmcm_locked(1);

      -- Input buffering
      --------------------------------------
    clkin1_buf : IBUFGDS
    port map (
        O  => clock_i,
        I  => clock_i_p,
        IB => clock_i_n
    );

    trigger_clocking : entity work.trigger_clocking
    port map(
        clk_in1           => clock_i,

        clk40_o           => clk_1x_gated_o,
        clk80_o           => clk_2x_gated_o,
        clk160_o          => clk_4x_gated_o,
        clk160_90_o       => clk_4x_90_gated_o,
        clk200_o          => clk_5x_gated_o,

        powerdown_i        => not clock_enable_i,

        locked_o          => mmcm_locked(0)
    );

    logic_clocking : entity work.logic_clocking
    port map(
        clk_in1     => clock_i,
        clk40_o     => clock,
        clk80_o     => clk_2x_o,
        clk160_0_o  => clk_4x_o,
        clk160_90_o => clk_4x_90_o,
        clk200_o    => clk_5x_o,
        locked_o    => mmcm_locked(1)
    );

    --===============================================================================================
    -- (this section is generated by <optohybrid_top>/tools/generate_registers.py -- do not edit)
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave_tmr
        generic map(
           g_NUM_REGS             => REG_CLOCKING_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_CLOCKING_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_CLOCKING_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => clock,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => clock,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_CLOCKING_ADDRESS_MSB downto REG_CLOCKING_ADDRESS_LSB) <= "00";

    -- Connect read signals
    regs_read_arr(0)(REG_CLOCKING_CORE_MMCM_LOCKED_BIT) <= mmcm_locked(1);
    regs_read_arr(0)(REG_CLOCKING_TRIGGER_MMCM_LOCKED_BIT) <= mmcm_locked(0);
    regs_read_arr(0)(REG_CLOCKING_CORE_MMCM_UNLOCKED_CNT_MSB downto REG_CLOCKING_CORE_MMCM_UNLOCKED_CNT_LSB) <= cnt_gbt_mmcm_unlocked;
    regs_read_arr(0)(REG_CLOCKING_TRIGGER_MMCM_UNLOCKED_CNT_MSB downto REG_CLOCKING_TRIGGER_MMCM_UNLOCKED_CNT_LSB) <= cnt_logic_mmcm_unlocked;

    -- Connect write signals

    -- Connect write pulse signals

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect counter instances

    COUNTER_CLOCKING_CORE_MMCM_UNLOCKED_CNT : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 8
    )
    port map (
        clk_i   => clock,
        rst_i   => ipb_reset_i,
        en_i    => mmcm_unlocked(1),
        snap_i  => '1',
        count_o => cnt_gbt_mmcm_unlocked
    );


    COUNTER_CLOCKING_TRIGGER_MMCM_UNLOCKED_CNT : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 8
    )
    port map (
        clk_i   => clock,
        rst_i   => ipb_reset_i,
        en_i    => mmcm_unlocked(0),
        snap_i  => '1',
        count_o => cnt_logic_mmcm_unlocked
    );


    -- Connect rate instances

    -- Connect read ready signals

    -- Defaults

    -- Define writable regs

    -- Create a sump for unused write signals
    sump_loop : for I in 0 to (REG_CLOCKING_NUM_REGS-1) generate
    begin
    regs_write_arr_sump (I) <= or_reduce (regs_write_arr(I));
    end generate;
    --==== Registers end ============================================================================

    --------------------------------------------------------------------------------------------------------------------
    -- Sump
    --------------------------------------------------------------------------------------------------------------------

    sump <= or_reduce(regs_write_arr_sump);

end Behavioral;
